float weight = 10.0;