sv name = "Marcelo";

function sayHello(name) {
    print("Hello");
    print("name");

    return 1;
}

sv expr = (10 * 10 + 10);

print("expr");
