switch(tk) {
    case "oi":
        print("OI");
        break;

    default:
        print("Hello");
}