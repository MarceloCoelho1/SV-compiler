switch(tk) {
    case "oi":
        print("OI");
        break;

    default:
        print("SALVE");
        break;
}


String name = "Marcelo";
char value = 'b';
int num = 10;
float num = 20.2;
bool name = true;


function sayHello(String name, int age) {
    print("Hello", name);
    print("Your age is: ", age);
}

sayHello("Marcelo", 19);