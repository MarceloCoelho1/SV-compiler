String name = "Marcelo";

function sayHello(name) {
    print("Hello");
    print(name);

    return 1;
}


int expr = (10 * 10 + 10);

print("expr");


if(true) {
    print("Hello");
} else {
    print("Hello");
}

while(true) {
    print("Hello");
    expr--;    
}

int name = 10;