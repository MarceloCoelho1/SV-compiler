switch(tk) {
    case "oi":
        print("OI");
        break;

    default:
        print("SALVE");
        break;
}


int value = (10 + 10 + 1);

String name = "Marcelo";
char value = 'b';
int num = 10;
float num = 20.2;
bool name = true;
double dsa = 20.1;

function sayHello(String name, int age) {
    print("Hello", name);
    print("Your age is: ", age);
}

sayHello("Marcelo", 19);

for (int i = 0; i < 10; i++) {
    print("oi");
}
