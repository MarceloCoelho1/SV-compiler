sv value = 10;